`define PRETRAINED
`define NUM_LAYERS 5
`define DATA_WIDTH 16
`define WEIGHT_INT_WIDTH 4
`define SIGMOID_SIZE 5

`define NUM_NEURON_L1 30
`define NUM_WEIGHT_L1 784
`define ACT_TYPE_L1 "relu"

`define NUM_NEURON_L2 30
`define NUM_WEIGHT_L2 30
`define ACT_TYPE_L2 "relu"

`define NUM_NEURON_L3 10
`define NUM_WEIGHT_L3 30
`define ACT_TYPE_L3 "relu"

`define NUM_NEURON_L4 10
`define NUM_WEIGHT_L4 10
`define ACT_TYPE_L4 "relu"

`define NUM_NEURON_L5 10
`define NUM_WEIGHT_L5 10
`define ACT_TYPE_L5 "hardmax"